`define CONSOLE_138K

